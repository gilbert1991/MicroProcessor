--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package SingleCycle_PKG is

TYPE DATA_MEMORY is ARRAY(0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
TYPE INSTRUCTION_MEMORY is ARRAY(0 TO 255) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
TYPE GENERAL_PURPOSE_REGISTER is ARRAY(0 TO 31) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
TYPE ALU_OPERATION is (O_ADD, O_SUB, O_AND, O_OR, O_NOR, O_SHL, O_SHR,O_BLT, O_BEQ, O_BNE, O_NULL);

-- type <new_type> is
--  record
--    <type_name>        : std_logic_vector( 7 downto 0);
--    <type_name>        : std_logic;
-- end record;
--
-- Declare constants
--
-- constant <constant_name>		: time := <time_unit> ns;
-- constant <constant_name>		: integer := <value;
--
-- Declare functions and procedure
--
-- function <function_name>  (signal <signal_name> : in <type_declaration>) return <type_declaration>;
-- procedure <procedure_name> (<type_declaration> <constant_name>	: in <type_declaration>);
--

end SingleCycle_PKG;

package body SingleCycle_PKG is

---- Example 1
--  function <function_name>  (signal <signal_name> : in <type_declaration>  ) return <type_declaration> is
--    variable <variable_name>     : <type_declaration>;
--  begin
--    <variable_name> := <signal_name> xor <signal_name>;
--    return <variable_name>; 
--  end <function_name>;

---- Example 2
--  function <function_name>  (signal <signal_name> : in <type_declaration>;
--                         signal <signal_name>   : in <type_declaration>  ) return <type_declaration> is
--  begin
--    if (<signal_name> = '1') then
--      return <signal_name>;
--    else
--      return 'Z';
--    end if;
--  end <function_name>;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;
 
end SingleCycle_PKG;
